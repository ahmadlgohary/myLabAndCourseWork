library verilog;
use verilog.vl_types.all;
entity circuit2_vlg_vec_tst is
end circuit2_vlg_vec_tst;
