library verilog;
use verilog.vl_types.all;
entity lab5circuit_vlg_vec_tst is
end lab5circuit_vlg_vec_tst;
