library verilog;
use verilog.vl_types.all;
entity CiruitProblem1_vlg_vec_tst is
end CiruitProblem1_vlg_vec_tst;
