library verilog;
use verilog.vl_types.all;
entity CiruitProblem3_vlg_vec_tst is
end CiruitProblem3_vlg_vec_tst;
