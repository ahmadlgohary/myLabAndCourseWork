library verilog;
use verilog.vl_types.all;
entity circuit_vlg_vec_tst is
end circuit_vlg_vec_tst;
